strict table
Unlimited stringtab-separated intI1-t-Required currencyC 2 USD1-1Up to 2 relative datesE-2
ValidRow1	212.345 3 BHDw+4.5
Tooshort
Toolong6	9	4204.20t+3h-1:23extra	field (1)extra field2
Wrongseparator89100.00
Missingrequiredvalueh-3
Incorrectcurrency8.8
another strict table
just one column this time
testrowwithmanyvalues
STRICT TABLE
testingthe return2

People who have a lot can afford to gamble.

People who have a little can’t afford to gamble.

People who have nothing can’t afford not to gamble. 

People who have a lot can afford to gamble.

People who have a little can’t afford to gamble.

People who have nothing can’t afford not to gamble. 
